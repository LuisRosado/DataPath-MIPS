module AND(
	input Din,Din2,
	output Dout
    );
	 
assign Dout = Din&Din2;

endmodule

